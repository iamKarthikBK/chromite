
/*
See LICENSE for details
This file has been generated by CSR-BOX - 1.5.4
Time of Generation: 2021-10-02 15:34:55.376148
*/

package csrbox;
   
import Vector           :: *;
import FIFOF            :: * ;
import DReg             :: * ;
import UniqueWrappers   :: * ;
import ConcatReg        :: * ;
import GetPut           :: * ;
import Connectable      :: * ;
import csr_types        :: * ;
import Assert           :: * ;
`include "csrbox.defines"
`include "Logger.bsv"
import csrbox_grp1 :: * ;
import csrbox_decoder :: * ;
  interface Sbread;
    method Bit#(64) mv_csr_misa;
    method Bit#(64) mv_csr_mvendorid;
    method Bit#(64) mv_csr_stvec;
    method Bit#(64) mv_csr_mtvec;
    method Bit#(64) mv_csr_mstatus;
    method Bit#(64) mv_csr_marchid;
    method Bit#(64) mv_csr_mimpid;
    method Bit#(64) mv_csr_mhartid;
    method Bit#(64) mv_csr_mip;
    method Bit#(64) mv_csr_sip;
    method Bit#(64) mv_csr_mie;
    method Bit#(64) mv_csr_sie;
    method Bit#(64) mv_csr_mscratch;
    method Bit#(64) mv_csr_sscratch;
    method Bit#(64) mv_csr_sepc;
    method Bit#(64) mv_csr_stval;
    method Bit#(64) mv_csr_scause;
    method Bit#(64) mv_csr_mepc;
    method Bit#(64) mv_csr_mtval;
    method Bit#(64) mv_csr_mcause;
    method Bit#(64) mv_csr_mcycle;
    method Bit#(64) mv_csr_minstret;
    method Bit#(64) mv_csr_time;
    method Bit#(64) mv_csr_mideleg;
    method Bit#(64) mv_csr_medeleg;
    method Bit#(64) mv_csr_pmpcfg0;
    method Bit#(64) mv_csr_pmpaddr0;
    method Bit#(64) mv_csr_pmpaddr1;
    method Bit#(64) mv_csr_pmpaddr2;
    method Bit#(64) mv_csr_pmpaddr3;
    method Bit#(64) mv_csr_satp;
    method Bit#(32) mv_csr_mcountinhibit;
    method Bit#(64) mv_csr_customcontrol;  
  endinterface:Sbread
  // Interaface declaration
  interface Ifc_csrbox;
    interface Sbread sbread;
    method Action ma_stop_count(Bit#(1) _stop);

    method Vector#(4, Bit#(8)) mv_pmpcfg;
    method Vector#(4, Bit#(32)) mv_pmpaddr;
    method Action ma_set_mip_meip (Bit#(1) _meip);
    method Action ma_set_mip_mtip (Bit#(1) _mtip);
    method Action ma_set_mip_msip (Bit#(1) _msip);
    method Action ma_set_mip_seip (Bit#(1) _seip);
    method Action ma_incr_minstret(Bit#(64) incr);
    method Action ma_set_time (Bit#(64) _time);
    method Action ma_set_mip_debug_interrupt (Bit#(1) _debug_interrupt);
    
    /*doc:method : to receive the request from the core or previous node" */
    method Action ma_core_req(CSRReq req); 

    /*doc:method : to send response to core on a hit in this node" */
    method CSRResponse mv_core_resp;

    method ActionValue#(Bit#(64)) mav_upd_on_ret (Bit#(8) retype);
    
    method ActionValue#(Bit#(64)) mav_upd_on_trap(Bit#(`causesize) cause, Bit#(64) pc, Bit#(64) tval);

    method Privilege_mode mv_prv;


  endinterface

  //Module Declarations
`ifdef csrbox_noinline
  (*synthesize*)
  
  (*conflict_free="ma_core_req,mv_core_resp"*)
(*conflict_free="ma_incr_minstret,sbread.mv_csr_minstret"*)
`endif
  module mk_csrbox(Ifc_csrbox);

    let grp1 <- mk_csrbox_grp1;

    let lv_misa_s = grp1.mv_csr_misa[18];
    let lv_misa_u = grp1.mv_csr_misa[20];
    let lv_misa_n = grp1.mv_csr_misa[13];
    let lv_misa_c = grp1.mv_csr_misa[2];
    /*doc:reg: holds the current privilege level*/
    Reg#(Privilege_mode) rg_prv <- mkReg(Machine);

    Bool anyhit = grp1.mv_core_resp.hit;
    Bit#(64) anydata = grp1.mv_core_resp.data;
    Wire#(Bit#(1)) wr_stop_count <- mkDWire(0);
    mkConnection(grp1.ma_stop_count, wr_stop_count);

    mkConnection(grp1.ma_upd_privilege, rg_prv);
    method ma_core_req = grp1.ma_core_req;
    method mv_core_resp = CSRResponse{hit:anyhit, data: anydata};
    method mv_prv = rg_prv;
    method ActionValue#(Bit#(64)) mav_upd_on_ret (Bit#(8) retype);
      Privilege_mode prv = unpack(retype[5:4]);
      Bool dret = (retype[3:0] == 'hb);
      Bit#(TSub#(64,1)) lv_epc = ?;

      if (prv == Supervisor) begin
        grp1.ma_set_mstatus_spie(1'b1);
        grp1.ma_set_mstatus_sie(grp1.mv_csr_mstatus[5]);
        rg_prv <= unpack(zeroExtend(grp1.mv_csr_mstatus[8]));
        lv_epc = truncateLSB(grp1.mv_csr_sepc);
        if (lv_misa_u == 1)
          grp1.ma_set_mstatus_spp(0);
        else
          grp1.ma_set_mstatus_spp(1);
        grp1.ma_set_mstatus_mprv(0);
      end
      else

      if (prv == Machine) begin
        grp1.ma_set_mstatus_mpie(1'b1);
        grp1.ma_set_mstatus_mie(grp1.mv_csr_mstatus[7]);
        rg_prv <= unpack(grp1.mv_csr_mstatus[12:11]);
        lv_epc = truncateLSB(grp1.mv_csr_mepc);
        if (lv_misa_u == 1)
          grp1.ma_set_mstatus_mpp(pack(User));
        else
          grp1.ma_set_mstatus_mpp(pack(Machine));
        if (grp1.mv_csr_mstatus[12:11] != '1)
          grp1.ma_set_mstatus_mprv(0);
      end
      if (lv_misa_c == 0)
        lv_epc[0] = 0;
      return {lv_epc, 1'b0};
    endmethod
    
    method ActionValue#(Bit#(64)) mav_upd_on_trap(Bit#(`causesize) cause, Bit#(64) pc, Bit#(64) tval);
      Bit#(TSub#(`causesize,1)) lv_cause = truncate(cause);
      Bit#(1) lv_trap_type = truncateLSB(cause);
      Bit#(64) lv_tvec = ?;
      Privilege_mode prv = Machine;
      Bool delegateM = False;
      Bool delegateS = False;

      let medeleg = grp1.mv_csr_medeleg;
      let mideleg = grp1.mv_csr_mideleg;
      delegateM = (truncate(mideleg >> lv_cause) & lv_trap_type) == 1 ||
                       (truncate(medeleg >> lv_cause) & ~lv_trap_type) == 1;

      if (delegateM && (pack(rg_prv) <= pack(Supervisor)) && (lv_misa_s == 1))
        prv = Supervisor;
      else if (delegateM && delegateS && rg_prv == User && lv_misa_n == 1 && lv_misa_s == 1)
        prv = User;
      else if (delegateM && rg_prv == User && lv_misa_n == 1 && lv_misa_s == 0)
        prv = User;

      if (prv == Supervisor) begin
        rg_prv <= Supervisor;
        grp1.ma_set_stval(tval);
        grp1.ma_set_sepc(pc);
        grp1.ma_set_scause({lv_trap_type, 'd0, lv_cause});
        grp1.ma_set_mstatus_sie(1'b0);
        grp1.ma_set_mstatus_spp(truncate(pack(rg_prv)));
        grp1.ma_set_mstatus_spie(grp1.mv_csr_mstatus[1]);
        Bit#(2) lv_trapmode = truncate(grp1.mv_csr_stvec);
        lv_tvec = {truncateLSB(grp1.mv_csr_stvec),2'b0};
        if ( lv_trapmode == 1 && lv_trap_type == 1)
          lv_tvec =  lv_tvec + {zeroExtend(lv_cause),2'b0};
      end
      else

      if (prv == Machine) begin
        rg_prv <= Machine;
        grp1.ma_set_mtval(tval);
        grp1.ma_set_mepc(pc);
        grp1.ma_set_mcause({lv_trap_type, 'd0, lv_cause});
        grp1.ma_set_mstatus_mie(1'b0);
        grp1.ma_set_mstatus_mpp(pack(rg_prv));
        grp1.ma_set_mstatus_mpie(grp1.mv_csr_mstatus[3]);
        Bit#(2) lv_trapmode = truncate(grp1.mv_csr_mtvec);
        lv_tvec = {truncateLSB(grp1.mv_csr_mtvec),2'b0};
        if ( lv_trapmode == 1 && lv_trap_type == 1)
            lv_tvec =  lv_tvec + {zeroExtend(lv_cause),2'b0};
      end
      return lv_tvec;
    endmethod
    method Action ma_stop_count(Bit#(1) _stop);
      wr_stop_count <= _stop;
    endmethod

    method Vector#(4, Bit#(32)) mv_pmpaddr;
        Vector#(4, Bit#(32)) lv_pmpaddr;
        lv_pmpaddr[0] = {truncate(grp1.mv_csr_pmpaddr0),2'b0};
        lv_pmpaddr[1] = {truncate(grp1.mv_csr_pmpaddr1),2'b0};
        lv_pmpaddr[2] = {truncate(grp1.mv_csr_pmpaddr2),2'b0};
        lv_pmpaddr[3] = {truncate(grp1.mv_csr_pmpaddr3),2'b0};

        return lv_pmpaddr;
    endmethod:mv_pmpaddr

    method Vector#(4, Bit#(8)) mv_pmpcfg;
        Vector#(4, Bit#(8)) lv_pmpcfg;
        lv_pmpcfg[0] = grp1.mv_csr_pmpcfg0[7:0];
        lv_pmpcfg[1] = grp1.mv_csr_pmpcfg0[15:8];
        lv_pmpcfg[2] = grp1.mv_csr_pmpcfg0[23:16];
        lv_pmpcfg[3] = grp1.mv_csr_pmpcfg0[31:24];

        return lv_pmpcfg;
    endmethod:mv_pmpcfg

    interface Sbread sbread;
      method mv_csr_misa = grp1.mv_csr_misa;

      method mv_csr_mvendorid = grp1.mv_csr_mvendorid;

      method mv_csr_stvec = grp1.mv_csr_stvec;

      method mv_csr_mtvec = grp1.mv_csr_mtvec;

      method mv_csr_mstatus = grp1.mv_csr_mstatus;

      method mv_csr_marchid = grp1.mv_csr_marchid;

      method mv_csr_mimpid = grp1.mv_csr_mimpid;

      method mv_csr_mhartid = grp1.mv_csr_mhartid;

      method mv_csr_mip = grp1.mv_csr_mip;

      method mv_csr_sip = grp1.mv_csr_sip;

      method mv_csr_mie = grp1.mv_csr_mie;

      method mv_csr_sie = grp1.mv_csr_sie;

      method mv_csr_mscratch = grp1.mv_csr_mscratch;

      method mv_csr_sscratch = grp1.mv_csr_sscratch;

      method mv_csr_sepc = grp1.mv_csr_sepc;

      method mv_csr_stval = grp1.mv_csr_stval;

      method mv_csr_scause = grp1.mv_csr_scause;

      method mv_csr_mepc = grp1.mv_csr_mepc;

      method mv_csr_mtval = grp1.mv_csr_mtval;

      method mv_csr_mcause = grp1.mv_csr_mcause;

      method mv_csr_mcycle = grp1.mv_csr_mcycle;

      method mv_csr_minstret = grp1.mv_csr_minstret;

      method mv_csr_time = grp1.mv_csr_time;

      method mv_csr_mideleg = grp1.mv_csr_mideleg;

      method mv_csr_medeleg = grp1.mv_csr_medeleg;

      method mv_csr_pmpcfg0 = grp1.mv_csr_pmpcfg0;

      method mv_csr_pmpaddr0 = grp1.mv_csr_pmpaddr0;

      method mv_csr_pmpaddr1 = grp1.mv_csr_pmpaddr1;

      method mv_csr_pmpaddr2 = grp1.mv_csr_pmpaddr2;

      method mv_csr_pmpaddr3 = grp1.mv_csr_pmpaddr3;

      method mv_csr_satp = grp1.mv_csr_satp;

      method mv_csr_mcountinhibit = grp1.mv_csr_mcountinhibit;

      method mv_csr_customcontrol = grp1.mv_csr_customcontrol;

    endinterface
    method ma_set_mip_meip = grp1.ma_set_mip_meip;
    method ma_set_mip_mtip = grp1.ma_set_mip_mtip;
    method ma_set_mip_msip = grp1.ma_set_mip_msip;
    method ma_set_mip_seip = grp1.ma_set_mip_seip;
    method ma_incr_minstret = grp1.ma_incr_minstret;
    method ma_set_time = grp1.ma_set_time;
    method ma_set_mip_debug_interrupt = grp1.ma_set_mip_debug_interrupt;
  endmodule 
endpackage 
