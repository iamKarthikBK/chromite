/*
Copyright (c) 2018, IIT Madras All rights reserved.

Redistribution and use in source and binary forms, with or without modification, are permitted
provided that the following conditions are met:

* Redistributions of source code must retain the above copyright notice, this list of conditions
  and the following disclaimer.  
* Redistributions in binary form must reproduce the above copyright notice, this list of 
  conditions and the following disclaimer in the documentation and/or other materials provided 
 with the distribution.  
* Neither the name of IIT Madras  nor the names of its contributors may be used to endorse or 
  promote products derived from this software without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS
OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER
IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT 
OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--------------------------------------------------------------------------------------------------
Author: Neel Gala,Deepa N. Sarma
Email id: neelgala@gmail.com
Details:
--------------------------------------------------------------------------------------------------
*/

package icache_dm;
  import icache_types::*;
  import mem_config::*;
  import GetPut::*;
  import FIFOF::*;
  import BUtils ::*;  
  import DReg::*;
  
  //parameters:
  // wordsize: number of bytes per word. This is what is responded back to the core.
  // blocksize: number of words per data line.
  // sets: number of sets within the cache.
  
  interface Ifc_icache_dm#(numeric type wordsize, numeric type blocksize,  numeric type sets,numeric
  type respwidth, numeric type paddr);
  interface Put#(ICore_request#(paddr)) core_req;
  interface Get#(ICore_response#(respwidth)) core_resp;
  interface Get#(IMem_request#(paddr)) mem_req;
  interface Put#(IMem_response#(respwidth)) mem_resp;
  `ifdef simulate
    interface Get#(Bit#(1)) meta;
  `endif
  endinterface

  (*conflict_free="check_hit_or_miss,poll_on_lb"*)
  (*preempts="get_io_response, check_hit_or_miss"*)
  module mkicache_dm#(function Bool is_IO(Bit#(paddr) addr))(Ifc_icache_dm#(wordsize,blocksize,sets,respwidth, paddr))
  provisos(
            Mul#(wordsize, 8, _w),        // _w is the total bits in a word
            Mul#(blocksize, _w,linewidth),// linewidth is the total bits in a cache line
            Log#(wordsize,wordbits),      // wordbits is no. of bits to index a byte in a word
            Log#(blocksize, blockbits),   // blockbits is no. of bits to index a word in a block
            Log#(sets, setbits),          // setbits is the no. of bits used as index in BRAMs.
            Add#(wordbits,blockbits,_a),  // _a total bits to index a byte in a cache line.
            Add#(_a, setbits, _b),        // _b total bits for index+offset, 
            Add#(tagbits, _b, paddr),        // tagbits = 32-(wordbits+blockbits+setbits)
            Mul#(wordsize,8,word_len),    // word_len = number of bits in a word
            Div#(respwidth,word_len,num_words),//num_words=number of words fetched from memory in a
            //cycle
            // Provisos for mem_config. If the number of banks have changed then the following
            // provisos will have to be re-written.
            Add#(a__, TDiv#(linewidth, 8), linewidth),
            Mul#(TDiv#(TDiv#(linewidth, 8), TDiv#(TDiv#(linewidth, 8), 8)),
              TDiv#(TDiv#(linewidth, 8), 8), TDiv#(linewidth, 8)),
            Mul#(TDiv#(linewidth, 8), 8, linewidth),
            // following provisos required by compiler:
            Bits#(Tuple2#(Bit#(respwidth), Bool), c__),
            Add#(d__, 1, blocksize),
            Add#(e__, respwidth, linewidth),
            Mul#(respwidth, f__, linewidth)
            );
  
    let v_sets=valueOf(sets);
    let v_setbits=valueOf(setbits);
    let v_wordbits=valueOf(wordbits);
    let v_blockbits=valueOf(blockbits);
    let v_linewidth=valueOf(linewidth);
    let v_tagbits=valueOf(tagbits);
    let v_num_words=valueOf(num_words);
    let verbosity=`VERBOSITY;
    let v_paddr=valueOf(paddr);
//    let paddr    = valueOf(PADDR);

    //Following function returns the info regarding word_position in line getting filled
    function Bit#(blocksize) fn_enable(Bit#(blockbits)word_index);
       Bit#(blocksize) write_enable ='h0; //
       for(Integer i=0;i<v_num_words;i=i+1)
         write_enable[word_index+fromInteger(i)]=1;
       return write_enable;
    endfunction

    Ifc_mem_config#(sets, linewidth, 8) data_arr <- mkmem_config_h; // data array
    Ifc_mem_config#(sets, TAdd#(1, tagbits), 1) tag_arr <- mkmem_config_h; // one extra valid bit
    
    FIFOF#(ICore_response#(respwidth))ff_core_response <- mkSizedFIFOF(2);
    FIFOF#(IMem_request#(paddr)) ff_mem_request    <- mkSizedFIFOF(2);
    FIFOF#(IMem_response#(respwidth)) ff_mem_response  <- mkSizedFIFOF(2);

    FIFOF#(ICore_request#(paddr)) ff_req_queue <- mkSizedFIFOF(2); 
    // The following fifo indicates if there is a miss that is pending a response to the core.
    FIFOF#(Bit#(paddr)) ff_miss_ongoing <- mkSizedFIFOF(1);
    FIFOF#(ICore_response#(respwidth)) ff_delayed_resp <- mkSizedFIFOF(1);

    `ifdef simulate
      FIFOF#(Bit#(1)) ff_meta <- mkSizedFIFOF(2);
      FIFOF#(Bit#(1)) ff_delayed_meta <- mkSizedFIFOF(1);
    `endif

    Reg#(Bit#(TLog#(sets))) rg_fence_index <- mkReg(0);
    Reg#(Bool) rg_init <- mkReg(True);
    Reg#(Bool) rg_fence_stall <- mkReg(True);
    Reg#(Bit#(blocksize))rg_blockenable <- mkReg(0);
    Reg#(Bit#(blockbits))index<-mkReg(0);
    //linebuffer control
    FIFOF#(Tuple3#(Bit#(tagbits), Bit#(setbits),Bit#(blocksize))) ff_lb_control <- mkUGSizedFIFOF(2);
    Reg#(Tuple4#(Bit#(1), Bit#(linewidth), Bit#(blocksize), Bool)) rg_linebuff <- 
                                                                      mkReg(tuple4(0, 0, 0, False));
    Reg#(Bool) rg_deq_lb <- mkDReg(False);

   
    // on reset we issue a fence instruction to initiliase the cache.
    rule initialize(rg_init);
      ff_req_queue.enq(tuple3(?,True,?));
      rg_init<=False;
    endrule


    //Fencing the cache
    // rule to fire only when there is not a pending fill to LB.
    // If this condition is not added then it is possible that LB populates the CACHE line after
    // being fenced which is wrong behavior
    rule fence_cache(tpl_2(ff_req_queue.first) && !ff_lb_control.notEmpty && rg_fence_stall);
       tag_arr.write_request(rg_fence_index,'d0);
       rg_fence_index<= rg_fence_index+1;
       if(verbosity>0)
         $display($time,"\tICACHE: Fence in progress. Index: %d",rg_fence_index);
       if(rg_fence_index==(fromInteger(v_sets-1))) begin
          ff_req_queue.deq;
          rg_fence_stall<=False;
          if(verbosity>1)begin
            $display($time,"\tICACHE Params:");
            $display($time,"\tv_sets: %d",v_sets);
            $display($time,"\tv_setbits: %d",v_setbits);
            $display($time,"\tv_wordbits: %d",v_wordbits);
            $display($time,"\tv_blockbits: %d",v_blockbits);
            $display($time,"\tv_tagbits: %d",v_tagbits);
            $display($time,"\tv_num_words: %d",v_num_words);
          end
       end
    endrule
    
    //Checking_line_buffer and cache
    rule check_hit_or_miss(!ff_delayed_resp.notEmpty && !tpl_2(ff_req_queue.first));
      //TODO: Should epochs be checked here also?
      let {request, fence, epoch} =ff_req_queue.first();
      ff_req_queue.deq;
      Bit#(TAdd#(3,TAdd#(wordbits,blockbits)))block_offset=
                                                          (request[v_blockbits+v_wordbits-1:0])<<3;
      Bit#(blockbits) word_index=request[v_blockbits+v_wordbits-1:v_wordbits];
      Bit#(linewidth) dataline <- data_arr.read_response;
      Bit#(TAdd#(1, tagbits)) tag <- tag_arr.read_response;
      Bit#(tagbits) request_tag = request[v_paddr-1:v_paddr-v_tagbits];
      Bit#(1) valid=tag[v_tagbits];
      Bit#(tagbits) stored_tag=tag[v_tagbits-1:0];
      let set_index=request[v_setbits+v_blockbits+v_wordbits-1:v_blockbits+v_wordbits];

      if(verbosity!=0)begin
        $display($time,"\tICACHE: Check for Address:%h Valid: %b ReqTag: %h StoredTag: %h",
            request,valid,request_tag,stored_tag);
      end

      let {lbvalid, lbdataline,lbenables,err} = rg_linebuff;
      let {lbtag,lbset,init_we}=ff_lb_control.first();

      // We first check if the requested word is in the line-buffer. This is done by checking the
      // if the tags match. While this means that the line-buffer should have the data
      // required, it might not be available unless it has been filled by the memory. We can confirm
      // this by checking the byte-enables which indicate which bytes of the line are available and
      // also confirm if the valid bit is set.

      // TODO check for IO request here before anything else.
      if(is_IO(request))begin
        if(verbosity>0)
          $display($time,"\tICACHE: This address is IO Mapped. Sending to memory");
        ff_mem_request.enq(tuple3(request,0,2));
        ff_miss_ongoing.enq(1);
      end
      else begin
        if(lbtag==request_tag && lbset==set_index && ff_lb_control.notEmpty) begin // hit in line-buffer
          if(verbosity!=0)
            $display($time,"\tICACHE: LB Holds the line for address: %h",request);
          if(lbenables[word_index]!=1||lbvalid!=1) begin
            if(verbosity!=0)
              $display($time,"\tICACHE: Miss. Word not found in LB for address: %h",request);
            ff_miss_ongoing.enq(request);
          end  
          else begin
            if(verbosity!=0)
              $display($time,"\tICACHE: Hit. Word present in LB");
            Bit#(respwidth) word_response = truncate(lbdataline>>block_offset); 

            if(ff_miss_ongoing.notEmpty) begin
              ff_delayed_resp.enq(tuple2(word_response,False));
              `ifdef simulate
                ff_delayed_meta.enq(1);
              `endif
            end
            else begin
              ff_core_response.enq(tuple2(word_response, False));// word and no bus-error;
              `ifdef simulate
                ff_meta.enq(1);
              `endif
            end
            if(verbosity!=0)
              $display($time,"\tICACHE: Sending the response back to the core from address:%h data:%h",
                request,word_response);
          end
        end
        else begin // since LB doesn't hold the required line check the cache.
          if((valid==1) && (stored_tag==request_tag)) begin // hit in cache
            Bit#(respwidth) word_response = truncate(dataline>>block_offset); 
            if(ff_miss_ongoing.notEmpty)begin
              ff_delayed_resp.enq(tuple2(word_response,False));
              `ifdef simulate
                ff_delayed_meta.enq(1);
              `endif
            end
            else begin
              ff_core_response.enq(tuple2(word_response, False));// word and no bus-error;
              `ifdef simulate
                ff_meta.enq(1);
              `endif
            end
            if(verbosity!=0)
              $display($time,"\tHIT IN CACHE for addr:%h data:%h",request,word_response);
          end
          else begin
            if(verbosity!=0)
                $display($time,"\tICACHE: Miss in Cache for addr: %h",request);
            ff_miss_ongoing.enq(request);
            ff_mem_request.enq(tuple3(request,fromInteger(valueOf(blocksize)-1),2));
            // TODO check if the following is valid.
            // Here we do not check if the lb_control is full since ff_req is of the same size and has
            // implicit condition on the rule. Thus if ff_req_queue is full then lb_control is also
            // full.
            ff_lb_control.enq(tuple3(request_tag,set_index,fn_enable(word_index)));
          end
        end        
      end
    endrule

    rule deque_delayed_response(!ff_miss_ongoing.notEmpty && ff_delayed_resp.notEmpty);
      if(verbosity>0)
        $display($time,"\tICACHE: Sending delayed response");
      ff_core_response.enq(ff_delayed_resp.first());
      ff_delayed_resp.deq;
      `ifdef simulate
        ff_meta.enq(ff_delayed_meta.first());
        ff_delayed_meta.deq;
      `endif
    endrule

    rule poll_on_lb(ff_lb_control.notEmpty);
      let {lbvalid, lbdataline,lbenables,err} = rg_linebuff;
      let {lbtag,lbset,init_we}=ff_lb_control.first();
      let request=ff_miss_ongoing.first();
      Bit#(tagbits) request_tag = request[v_paddr-1:v_paddr-v_tagbits]; 
      let set_index=request[v_setbits+v_blockbits+v_wordbits-1:v_blockbits+v_wordbits];
      Bit#(blockbits) word_index=request[v_blockbits+v_wordbits-1:v_wordbits];
      Bit#(TAdd#(3,TAdd#(wordbits,blockbits)))block_offset=
                                                          (request[v_blockbits+v_wordbits-1:0])<<3;

      if(lbtag==request_tag && lbset==set_index && ff_lb_control.notEmpty) begin // hit in line-buffer
        if(verbosity!=0)
          $display($time,"\tICACHE: Polling LB Holds the line for address: %h",request);
        if(lbenables[word_index]!=1||lbvalid!=1) begin
          if(verbosity!=0)
            $display($time,"\tICACHE: Polling Miss. Word not found in LB for address: %h",request);
        end  
        else begin
          if(verbosity!=0)
              $display($time,"\tICACHE: Polling Hit. Word present in LB for address: %h",request);
          Bit#(respwidth) word_response = truncate(lbdataline>>block_offset); 
          ff_core_response.enq(tuple2(word_response,err));// word and no bus-error;
          `ifdef simulate
            ff_meta.enq(0);
          `endif
          ff_miss_ongoing.deq;
          if(verbosity!=0)
            $display($time,"\tICACHE: Polling Sending the response back to the core from address:%h data:%h",
              request,word_response);
        end
      end
    endrule
    
    //Reading IO_response
    // TODO: When should this fire?
    rule get_io_response(!ff_lb_control.notEmpty);
      let {word,err} = ff_mem_response.first;
      if(verbosity>0)
        $display($time,"\tICACHE: receiving IO response: %h",word);
      ff_mem_response.deq;
      ff_core_response.enq(tuple2(word, err));// word and no bus-error;
      `ifdef simulate
        ff_meta.enq(0);
      `endif
      ff_miss_ongoing.deq();
    endrule

    //Capturing memory_response
    rule capture_memory_response(&(tpl_3(rg_linebuff))!=1 && ff_lb_control.notEmpty);
     
      Bit#(linewidth) mask = 0;
      let {word,err} = ff_mem_response.first;
      ff_mem_response.deq;
      if (verbosity!=0)
        $display($time,"\tICACHE: Receiving Memory Response. Word: %h err: %b",word,err);
      let {lbvalid, lbdataline,lbenables, err1} = rg_linebuff;
      let {lbtag,lbset, init_we}=ff_lb_control.first();
      Bit#(blocksize) temp = 0;
      if(rg_blockenable==0)
        temp=init_we;
      else
        temp=rg_blockenable;

      lbenables = lbenables|temp;

      if (verbosity!=0)
        $display($time,"\tICACHE: Lbenables changes to:%b",lbenables);

      rg_blockenable <= {temp[valueOf(blocksize)-2:0],
                                                temp[valueOf(blocksize)-1]};

      if (verbosity!=0)
        $display($time,"\tICACHE: WE :%b",temp);

     //Each bit in write_enable register refers to corresponding word in block 
      
      for(Integer i=0;i<valueOf(blocksize);i=i+1)
      begin
            Bit#(respwidth) ex_we=duplicate(temp[i]);
            let v_word_len = valueOf(word_len);
            mask[((i*v_word_len)+(v_word_len-1)):i*v_word_len]=ex_we;
      end

      if (verbosity!=0)
        $display($time,"\tICACHE: MASK:%h",mask);

      Bit#(linewidth) y  = duplicate(word) ; 
      let new_word_line  = y & mask;
      Bit#(linewidth) x  = lbdataline|new_word_line;
      rg_linebuff <= tuple4(1'b1,x,lbenables, err||err1);

      if(verbosity!=0)
        $display($time,"\tICACHE: Updating line_buffer:%h",x);

    endrule

    //Loading data into the cache from line_buffer
    rule upd_data_into_cache(&(tpl_3(rg_linebuff))==1 && (tpl_1(rg_linebuff)==1) &&
                                                  ff_lb_control.notEmpty  && !rg_deq_lb);

      let {lbtag,lbset,init_we}=ff_lb_control.first();
      tag_arr.write_request(lbset,{1,lbtag});//lbtag
      data_arr.write_request(lbset,truncate(tpl_2(rg_linebuff)));
      if(verbosity!=0)
        $display($time,"\tICACHE: loading set:%h with dataline %h and tag %h",
                                        lbset,tpl_2(rg_linebuff),lbtag);
      rg_deq_lb<=True;
    endrule
    rule deq_lb(rg_deq_lb && &(tpl_3(rg_linebuff))==1 && (tpl_1(rg_linebuff)==1) &&
                                                                        ff_lb_control.notEmpty);
      ff_lb_control.deq;
      rg_blockenable<=0;
      rg_linebuff<=tuple4(0,0,0, False);
    endrule

    interface core_req=interface Put
      method Action put(ICore_request#(paddr) req) if(!rg_init && !rg_fence_stall &&
      !ff_miss_ongoing.notEmpty);
        // TODO check if epochs match. If they do not then drop the request.
        let {addr, fence, epoch} =req;
        if(fence)
          rg_fence_stall<=True;
        if (verbosity!=0)
		    $display($time,"\tICACHE: Receiving request to address:%h Fence: %b epoch: %b ",addr, fence,
                  epoch); 

        ff_req_queue.enq(req);
        Bit#(setbits) set_index=addr[v_setbits+v_blockbits+v_wordbits-1:v_blockbits+v_wordbits];
        data_arr.read_request(set_index);
        tag_arr.read_request(set_index);
        if(verbosity!=0)
		      $display($time,"\tICACHE: Access Cache for Addr: %h Index: %d",addr,set_index); 
        
      endmethod
    endinterface;

    interface core_resp = interface Get
      method ActionValue#(ICore_response#(respwidth)) get();
        ff_core_response.deq;
        return ff_core_response.first;
      endmethod
    endinterface;
    
    interface mem_req = interface Get
      method ActionValue#(IMem_request#(paddr)) get;
        ff_mem_request.deq;
        return ff_mem_request.first;
      endmethod
    endinterface;

    interface mem_resp= interface Put
     method Action put(IMem_response#(respwidth) resp);
        ff_mem_response.enq(resp);
     endmethod
    endinterface;
    `ifdef simulate 
      interface meta = interface Get
        method ActionValue#(Bit#(1)) get();
          ff_meta.deq;
          return ff_meta.first;
        endmethod
      endinterface;
    `endif 

  endmodule

endpackage
