
/* 
Copyright (c) 2018, InCore Semiconductors All rights reserved.

Redistribution and use in source and binary forms, with or without modification, are permitted
provided that the following conditions are met:

* Redistributions of source code must retain the above copyright notice, this list of conditions
  and the following disclaimer.  
* Redistributions in binary form must reproduce the above copyright notice, this list of 
  conditions and the following disclaimer in the documentation and/or other materials provided 
 with the distribution.  
* Neither the name of InCore Semiconductors Pvt. Ltd.  nor the names of its contributors may be used to endorse or 
  promote products derived from this software without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS
OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY
AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER
IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT 
OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--------------------------------------------------------------------------------------------------

Author: Vishvesh Sundararaman
Email id: vishu.vivek@gmail.com
Details:

mmap-start
slave_bound: 128 bytes

schema-start
module:
    type: string
    regex: ^sdram$
type:
    type: string
    regex: ^device$
clusters:
    type: list
    schema:
        type: string
roles:
    type: dict
    schema:
        master:
            type: list
            schema:
                type: string
                regex: ^(null$
                nullable: True
        slave:
            type: list
parameters:
    type: dict
    schema:
        clock:
            type: integer
            min: 1
            max: 1
        io_width:
            type: integer
            max: 64
        rfrsh_timer_width:
            type: integer
        rfrsh_row_width:
            type: integer
schema-end
*/

package sdram_template;
import sdram::*;
`include "sdram.defines"
import device_common::*;

(*synthesize*)
module mkdummy#(Clock sdram_clock, Reset sdram_reset)(Empty);
	let core_clock<-exposeCurrentClock;
	let core_reset<-exposeCurrentReset;
	Ifc_sdram_axi4#(32,64,0,64,12,3) sdram <- mksdram_axi4(sdram_clock,sdram_reset);

    rule rl_ipad;
     sdram.io.ipad_sdr_din(?);
    endrule
endmodule

endpackage
    
